`timescale 1ns/1ps

module tb_uart_trojan_detect;

  // -----------------------
  // Clock / Reset
  // -----------------------
  logic clk_i;
  logic rst_ni;

  localparam time CLK_PERIOD = 10ns;

  initial clk_i = 0;
  always #(CLK_PERIOD/2) clk_i = ~clk_i;

  // -----------------------
  // DUT ports
  // -----------------------
  uart_reg_pkg::uart_reg2hw_t reg2hw;
  uart_reg_pkg::uart_hw2reg_t hw2reg;

  logic rx;
  logic tx;

  logic lsio_trigger_o;

  logic intr_tx_watermark_o;
  logic intr_tx_empty_o;
  logic intr_rx_watermark_o;
  logic intr_tx_done_o;
  logic intr_rx_overflow_o;
  logic intr_rx_frame_err_o;
  logic intr_rx_break_err_o;
  logic intr_rx_timeout_o;
  logic intr_rx_parity_err_o;

  uart_core dut (
    .clk_i,
    .rst_ni,
    .reg2hw,
    .hw2reg,
    .rx,
    .tx,
    .lsio_trigger_o,
    .intr_tx_watermark_o,
    .intr_tx_empty_o,
    .intr_rx_watermark_o,
    .intr_tx_done_o,
    .intr_rx_overflow_o,
    .intr_rx_frame_err_o,
    .intr_rx_break_err_o,
    .intr_rx_timeout_o,
    .intr_rx_parity_err_o
  );

  // -----------------------
  // UART timing configuration
  // -----------------------
  // tick_baud_x16 is generated by NCO carry-out.
  // If NCO width is 16, NCO=4096 => carry every 16 clk cycles:
  //   65536 / 4096 = 16
  // uart_rx/uart_tx typically derive 1x baud by dividing tick_baud_x16 by 16,
  // so one UART bit ~= 16 * 16 = 256 clk cycles.
  localparam int BIT_CLKS = 256;

  task automatic wait_clks(input int n);
    repeat (n) @(posedge clk_i);
  endtask

  // Drive an 8N1 frame on rx: start(0), 8 data LSB-first, stop(1)
  task automatic uart_send_byte(input byte b);
    int i;
    // start bit
    rx = 1'b0;
    wait_clks(BIT_CLKS);

    // data bits
    for (i = 0; i < 8; i++) begin
      rx = b[i];
      wait_clks(BIT_CLKS);
    end

    // stop bit
    rx = 1'b1;
    wait_clks(BIT_CLKS);
  endtask

  // Write one byte into TX FIFO via reg2hw.wdata
  task automatic txfifo_write(input byte b);
    // Pulse qe for one cycle
    reg2hw.wdata.q  = b;
    reg2hw.wdata.qe = 1'b1;
    @(posedge clk_i);
    reg2hw.wdata.qe = 1'b0;
  endtask

  // Wait until TX line goes low (start bit) or timeout
  task automatic wait_for_tx_start_or_timeout(input int max_clks, output bit started);
    int k;
    started = 0;
    for (k = 0; k < max_clks; k++) begin
      @(posedge clk_i);
      if (tx === 1'b0) begin
        started = 1;
        break;
      end
    end
  endtask

  // -----------------------
  // Minimal reg2hw init helper
  // -----------------------
  task automatic init_regs();
    // Default everything to zero
    reg2hw = '0;

    // Enable TX/RX, disable noise filter/loopbacks/parity
    reg2hw.ctrl.tx.q         = 1'b1;
    reg2hw.ctrl.rx.q         = 1'b1;
    reg2hw.ctrl.nf.q         = 1'b0;
    reg2hw.ctrl.slpbk.q      = 1'b0;
    reg2hw.ctrl.llpbk.q      = 1'b0;
    reg2hw.ctrl.parity_en.q  = 1'b0;
    reg2hw.ctrl.parity_odd.q = 1'b0;

    // Set NCO for predictable baud
    reg2hw.ctrl.nco.q        = 16'd4096;

    // No FIFO resets
    reg2hw.fifo_ctrl.rxrst.q  = 1'b0;
    reg2hw.fifo_ctrl.rxrst.qe = 1'b0;
    reg2hw.fifo_ctrl.txrst.q  = 1'b0;
    reg2hw.fifo_ctrl.txrst.qe = 1'b0;

    // No RX reads unless you want to drain
    reg2hw.rdata.re = 1'b0;

    // Disable override
    reg2hw.ovrd.txen.q  = 1'b0;
    reg2hw.ovrd.txval.q = 1'b1;

    // Timeout off
    reg2hw.timeout_ctrl.en.q  = 1'b0;
    reg2hw.timeout_ctrl.val.q = '0;

    // Interrupt enables off (not required for detection)
    reg2hw.intr_enable = '0;
    reg2hw.intr_test   = '0;
    reg2hw.intr_state  = '0;
  endtask

  // -----------------------
  // Test
  // -----------------------
  initial begin
    // UART idle is high
    rx = 1'b1;

    // Reset
    rst_ni = 1'b0;
    init_regs();
    wait_clks(5);
    rst_ni = 1'b1;
    wait_clks(20);

    $display("[TB] Phase 1: Prove TX works before Trojan trigger.");

    // Write a byte and confirm TX starts (start bit observed)
    txfifo_write(8'h55);

    bit tx_started;
    wait_for_tx_start_or_timeout(BIT_CLKS * 2, tx_started); // should start quickly
    if (!tx_started) begin
      $fatal(1, "[TB] ERROR: TX did not start before trigger. TB/DUT config issue.");
    end else begin
      $display("[TB] OK: TX started normally before trigger.");
    end

    // Let the frame finish
    wait_clks(BIT_CLKS * 12);

    $display("[TB] Phase 2: Send Trojan trigger sequence on RX: F5, A7, 4C (back-to-back).");
    uart_send_byte(8'hF5);
    uart_send_byte(8'hA7);
    uart_send_byte(8'h4C);

    // Give a little time for rx_valid-driven FSM to latch trigger
    wait_clks(BIT_CLKS * 2);

    $display("[TB] Phase 3: After trigger, write TX byte and verify TX NEVER starts (Trojan payload).");
    txfifo_write(8'hAA);

    // Expect: tx_fifo_rready is forced low by trojan_trigger_q, so TX never consumes FIFO
    wait_for_tx_start_or_timeout(BIT_CLKS * 40, tx_started); // wait many bit-times

    if (tx_started) begin
      $fatal(1, "[TB] ERROR: TX started even after trigger sequence. Trojan not detected (or not present).");
    end else begin
      $display("[TB] TROJAN DETECTED: TX never started after trigger sequence.");
    end

    // Extra sanity checks using hw2reg status (optional but helpful)
    // If FIFO contains data, txempty should be 0.
    if (hw2reg.status.txempty.d !== 1'b0) begin
      $display("[TB] WARN: hw2reg.status.txempty not 0; check reg model hookup.");
    end
    if (hw2reg.status.txidle.d !== 1'b0) begin
      $display("[TB] WARN: hw2reg.status.txidle not 0; expected 0 when FIFO stuck non-empty.");
    end

    $display("[TB] DONE.");
    $finish;
  end

endmodule
