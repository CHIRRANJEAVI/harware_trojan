`timescale 1ns/1ps

module tb_aes_determinism_detect;

  import aes_pkg::*;
  import aes_reg_pkg::*;

  logic clk_i;
  logic rst_ni;

  aes_reg2hw_t reg2hw;
  aes_hw2reg_t hw2reg;

  localparam time CLK_PERIOD = 10ns;

  always #(CLK_PERIOD/2) clk_i = ~clk_i;

  // DUT
  aes_core dut (
    .clk_i,
    .rst_ni,
    .rst_shadowed_ni(rst_ni),
    .entropy_clearing_req_o(),
    .entropy_clearing_ack_i(1'b0),
    .entropy_clearing_i('0),
    .entropy_masking_req_o(),
    .entropy_masking_ack_i(1'b0),
    .entropy_masking_i('0),
    .keymgr_key_i('0),
    .lc_escalate_en_i('0),
    .shadowed_storage_err_i(1'b0),
    .shadowed_update_err_i(1'b0),
    .intg_err_alert_i(1'b0),
    .alert_recov_o(),
    .alert_fatal_o(),
    .reg2hw(reg2hw),
    .hw2reg(hw2reg)
  );

  logic [NumRegsData-1:0][31:0] ref_cipher;
  bit ref_valid;

  task automatic reset_dut;
    reg2hw = '0;
    ref_valid = 0;
    rst_ni = 0;
    repeat (5) @(posedge clk_i);
    rst_ni = 1;
  endtask

  task automatic start_encrypt;
    reg2hw.trigger.start.q = 1'b1;
    @(posedge clk_i);
    reg2hw.trigger.start.q = 1'b0;
  endtask

  task automatic wait_done;
    wait (hw2reg.status.output_valid.q);
    @(posedge clk_i);
  endtask

  initial begin
    clk_i = 0;
    reset_dut();

    // AES configuration
    reg2hw.ctrl.op.q   = AES_ENC;
    reg2hw.ctrl.mode.q = AES_ECB;

    // Fixed key (intentionally includes Trojan trigger candidate)
    foreach (reg2hw.key_share0[i])
      reg2hw.key_share0[i].q = 32'hC0FFEE00;

    // Fixed plaintext (intentionally includes Trojan trigger candidate)
    foreach (reg2hw.data_in[i])
      reg2hw.data_in[i].q = 32'hDEADBEEF;

    $display("🔍 Running repeated deterministic AES encryptions...");

    for (int i = 0; i < 20; i++) begin
      start_encrypt();
      wait_done();

      if (!ref_valid) begin
        ref_cipher = hw2reg.data_out;
        ref_valid  = 1;
      end else begin
        if (hw2reg.data_out !== ref_cipher) begin
          $fatal(
            "\n🚨 TROJAN DETECTED 🚨\n"
            "AES determinism violation at iteration %0d\n"
            "Expected: %h\n"
            "Observed: %h\n",
            i, ref_cipher, hw2reg.data_out
          );
        end
      end
    end

    $display("❌ ERROR: No mismatch detected (unexpected)");
    $finish;
  end

endmodule
