// Stub testbench
// Extend to activate Trojan trigger
module tb;
initial begin
  #1000 $finish;
end
endmodule
